
`timescale 1 ns / 1 ps

module QEA_AXI #
(
	// Users to add parameters here
    parameter PE_NUM_WIDTH            = 2,
    parameter PE_NUM                  = 4,
    parameter DATA_WIDTH              = 32,
    parameter MAX_QBIT_WIDTH          = 6,
    parameter ALU_DATA_WIDTH          = DATA_WIDTH,
    parameter STATE_DATA_WIDTH        = DATA_WIDTH*2,
    parameter STATE_ADDR_WIDTH        = 16,
    parameter GATE_DATA_WIDTH         = DATA_WIDTH*2,
    parameter GATE_ADDR_WIDTH         = 6,
    parameter GATE_CONTEXT_DATA_WIDTH = DATA_WIDTH*2,
    parameter GATE_CONTEXT_ADDR_WIDTH = 6,
	parameter GATE_NUM_WIDTH          = 4,
	parameter NUM_FRAC_BIT            = 30,
	// parameter AXI_DATA_WIDTH		  = 256, 

	parameter START_BASE_PHYS  = 32'h08000000,
	parameter FINISH_BASE_PHYS = 32'h0C000000,
	parameter CTX_BASE_PHYS    = 32'h80000000,
	parameter STATE_BASE_PHYS  = 32'hC0000000,
	// User parameters ends
	// Do not modify the parameters beyond this line


	// Parameters of Axi Slave Bus Interface S00_AXI
	parameter integer C_S00_AXI_ID_WIDTH	= 1,
	parameter integer C_S00_AXI_DATA_WIDTH	= 256,
	parameter integer C_S00_AXI_ADDR_WIDTH	= 32,
	parameter integer C_S00_AXI_AWUSER_WIDTH	= 0,
	parameter integer C_S00_AXI_ARUSER_WIDTH	= 0,
	parameter integer C_S00_AXI_WUSER_WIDTH	= 0,
	parameter integer C_S00_AXI_RUSER_WIDTH	= 0,
	parameter integer C_S00_AXI_BUSER_WIDTH	= 0
)
(
	// Users to add ports here

	// User ports ends
	// Do not modify the ports beyond this line


	// Ports of Axi Slave Bus Interface S00_AXI
	input wire  s00_axi_aclk,
	input wire  s00_axi_aresetn,
	input wire [C_S00_AXI_ID_WIDTH-1 : 0] s00_axi_awid,
	input wire [C_S00_AXI_ADDR_WIDTH-1 : 0] s00_axi_awaddr,
	input wire [7 : 0] s00_axi_awlen,
	input wire [2 : 0] s00_axi_awsize,
	input wire [1 : 0] s00_axi_awburst,
	input wire  s00_axi_awlock,
	input wire [3 : 0] s00_axi_awcache,
	input wire [2 : 0] s00_axi_awprot,
	input wire [3 : 0] s00_axi_awqos,
	input wire [3 : 0] s00_axi_awregion,
	input wire [C_S00_AXI_AWUSER_WIDTH-1 : 0] s00_axi_awuser,
	input wire  s00_axi_awvalid,
	output wire  s00_axi_awready,
	input wire [C_S00_AXI_DATA_WIDTH-1 : 0] s00_axi_wdata,
	input wire [(C_S00_AXI_DATA_WIDTH/8)-1 : 0] s00_axi_wstrb,
	input wire  s00_axi_wlast,
	input wire [C_S00_AXI_WUSER_WIDTH-1 : 0] s00_axi_wuser,
	input wire  s00_axi_wvalid,
	output wire  s00_axi_wready,
	output wire [C_S00_AXI_ID_WIDTH-1 : 0] s00_axi_bid,
	output wire [1 : 0] s00_axi_bresp,
	output wire [C_S00_AXI_BUSER_WIDTH-1 : 0] s00_axi_buser,
	output wire  s00_axi_bvalid,
	input wire  s00_axi_bready,
	input wire [C_S00_AXI_ID_WIDTH-1 : 0] s00_axi_arid,
	input wire [C_S00_AXI_ADDR_WIDTH-1 : 0] s00_axi_araddr,
	input wire [7 : 0] s00_axi_arlen,
	input wire [2 : 0] s00_axi_arsize,
	input wire [1 : 0] s00_axi_arburst,
	input wire  s00_axi_arlock,
	input wire [3 : 0] s00_axi_arcache,
	input wire [2 : 0] s00_axi_arprot,
	input wire [3 : 0] s00_axi_arqos,
	input wire [3 : 0] s00_axi_arregion,
	input wire [C_S00_AXI_ARUSER_WIDTH-1 : 0] s00_axi_aruser,
	input wire  s00_axi_arvalid,
	output wire  s00_axi_arready,
	output wire [C_S00_AXI_ID_WIDTH-1 : 0] s00_axi_rid,
	output wire [C_S00_AXI_DATA_WIDTH-1 : 0] s00_axi_rdata,
	output wire [1 : 0] s00_axi_rresp,
	output wire  s00_axi_rlast,
	output wire [C_S00_AXI_RUSER_WIDTH-1 : 0] s00_axi_ruser,
	output wire  s00_axi_rvalid,
	input wire  s00_axi_rready
);
	// Instantiation of Axi Bus Interface S00_AXI
	AXI_Interface # ( 
        .PE_NUM_WIDTH(PE_NUM_WIDTH),
        .PE_NUM(PE_NUM),
        .DATA_WIDTH(DATA_WIDTH),
        .MAX_QBIT_WIDTH(MAX_QBIT_WIDTH),
        .ALU_DATA_WIDTH(ALU_DATA_WIDTH),
        .STATE_DATA_WIDTH(STATE_DATA_WIDTH),
        .STATE_ADDR_WIDTH(STATE_ADDR_WIDTH),
        .GATE_DATA_WIDTH(GATE_DATA_WIDTH),
        .GATE_ADDR_WIDTH(GATE_ADDR_WIDTH),
        .GATE_CONTEXT_DATA_WIDTH(GATE_CONTEXT_DATA_WIDTH),
        .GATE_CONTEXT_ADDR_WIDTH(GATE_CONTEXT_ADDR_WIDTH),
        .GATE_NUM_WIDTH(GATE_NUM_WIDTH),
        .NUM_FRAC_BIT(NUM_FRAC_BIT),
		.START_BASE_PHYS(START_BASE_PHYS),
		.FINISH_BASE_PHYS(FINISH_BASE_PHYS),
		.STATE_BASE_PHYS(STATE_BASE_PHYS),
		.CTX_BASE_PHYS(CTX_BASE_PHYS),

		.C_S_AXI_ID_WIDTH(C_S00_AXI_ID_WIDTH),
		.C_S_AXI_DATA_WIDTH(C_S00_AXI_DATA_WIDTH),
		.C_S_AXI_ADDR_WIDTH(C_S00_AXI_ADDR_WIDTH),
		.C_S_AXI_AWUSER_WIDTH(C_S00_AXI_AWUSER_WIDTH),
		.C_S_AXI_ARUSER_WIDTH(C_S00_AXI_ARUSER_WIDTH),
		.C_S_AXI_WUSER_WIDTH(C_S00_AXI_WUSER_WIDTH),
		.C_S_AXI_RUSER_WIDTH(C_S00_AXI_RUSER_WIDTH),
		.C_S_AXI_BUSER_WIDTH(C_S00_AXI_BUSER_WIDTH)
	) AXI_Interface (
		.S_AXI_ACLK(s00_axi_aclk),
		.S_AXI_ARESETN(s00_axi_aresetn),
		.S_AXI_AWID(s00_axi_awid),
		.S_AXI_AWADDR(s00_axi_awaddr),
		.S_AXI_AWLEN(s00_axi_awlen),
		.S_AXI_AWSIZE(s00_axi_awsize),
		.S_AXI_AWBURST(s00_axi_awburst),
		.S_AXI_AWLOCK(s00_axi_awlock),
		.S_AXI_AWCACHE(s00_axi_awcache),
		.S_AXI_AWPROT(s00_axi_awprot),
		.S_AXI_AWQOS(s00_axi_awqos),
		.S_AXI_AWREGION(s00_axi_awregion),
		.S_AXI_AWUSER(s00_axi_awuser),
		.S_AXI_AWVALID(s00_axi_awvalid),
		.S_AXI_AWREADY(s00_axi_awready),
		.S_AXI_WDATA(s00_axi_wdata),
		.S_AXI_WSTRB(s00_axi_wstrb),
		.S_AXI_WLAST(s00_axi_wlast),
		.S_AXI_WUSER(s00_axi_wuser),
		.S_AXI_WVALID(s00_axi_wvalid),
		.S_AXI_WREADY(s00_axi_wready),
		.S_AXI_BID(s00_axi_bid),
		.S_AXI_BRESP(s00_axi_bresp),
		.S_AXI_BUSER(s00_axi_buser),
		.S_AXI_BVALID(s00_axi_bvalid),
		.S_AXI_BREADY(s00_axi_bready),
		.S_AXI_ARID(s00_axi_arid),
		.S_AXI_ARADDR(s00_axi_araddr),
		.S_AXI_ARLEN(s00_axi_arlen),
		.S_AXI_ARSIZE(s00_axi_arsize),
		.S_AXI_ARBURST(s00_axi_arburst),
		.S_AXI_ARLOCK(s00_axi_arlock),
		.S_AXI_ARCACHE(s00_axi_arcache),
		.S_AXI_ARPROT(s00_axi_arprot),
		.S_AXI_ARQOS(s00_axi_arqos),
		.S_AXI_ARREGION(s00_axi_arregion),
		.S_AXI_ARUSER(s00_axi_aruser),
		.S_AXI_ARVALID(s00_axi_arvalid),
		.S_AXI_ARREADY(s00_axi_arready),
		.S_AXI_RID(s00_axi_rid),
		.S_AXI_RDATA(s00_axi_rdata),
		.S_AXI_RRESP(s00_axi_rresp),
		.S_AXI_RLAST(s00_axi_rlast),
		.S_AXI_RUSER(s00_axi_ruser),
		.S_AXI_RVALID(s00_axi_rvalid),
		.S_AXI_RREADY(s00_axi_rready)
	);

	// Add user logic here

	// User logic ends
endmodule
